module and_gate_gate_primitive (A, B, X);

  input A, B;
  output X;

  and U0(X, A, B);

endmodule
