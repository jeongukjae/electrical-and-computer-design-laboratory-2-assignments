module test(A, X);
  input A;
  output X;
  
  wire X;

  assign X = !A;

endmodule
